`timescale 1ns/10ps

// Test bench module
module tb_macc;

// Input Array
/////////////////////////////////////////////////////////
//                  Test Bench Signals                 //
/////////////////////////////////////////////////////////

reg clk;

/////////////////////////////////////////////////////////
//                  I/O Declarations                   //
/////////////////////////////////////////////////////////
// declare variables to hold signals going into submodule
reg signed [7:0] inA, inB;
reg macc_clear;

// Output Signals
wire signed [18:0] out;
reg [18:0]test_product;
reg [18:0]accumulate ;
integer i;

/////////////////////////////////////////////////////////
//              Submodule Instantiation                //
/////////////////////////////////////////////////////////

/*****************************************
RENAME SIGNALS TO MATCH YOUR MODULE
******************************************/
MAC DUT
(
    .clk        (clk),
    .macc_clear (macc_clear),
    .inA        (inA),
    .inB        (inB),
    .out    (out)
  );

initial begin
    // YOUR CODE GOES HERE
	 clk = 0;
	 inA = 8'b01111111;
	 inB = 8'b01111111;
	  
	 accumulate = 0;
	 
	 for(i = 0; i <= 2; i = i + 1) begin
	 test_product = inA * inB;
	 accumulate = accumulate + test_product;
	 end 
	 macc_clear = 1'b1;
	 #20
	 macc_clear = 1'b0;
	 #300
//Finish test with 127 * 127
//Start test with -128 * 127
	 
 	 inA = 8'b10000000;
	 inB = 8'b01111111;
	 accumulate = 0;
	 for(i = 0; i <= 1; i = i + 1) begin
	 test_product = inA * inB;
	 accumulate = accumulate + test_product;
	 end 
	 macc_clear = 1'b1;
	 #20
	macc_clear = 1'b0;
	#300
//Finish test with -128 * 127
//Start random case tests 
	for(i = 0; i <= 9; i = i + 1) begin
	inA = $random;
	inB = $random;
	accumulate = 0;
	test_product = inA * inB;
	accumulate = accumulate + test_product;
	#20
	macc_clear = 1'b1;
	#40
	macc_clear = 1'b0;
	
 	end
	 
	
	 
	
		
    $stop; // End Simulation

end

// Clock
always begin
   #10;           // wait for initial block to initialize clock
   clk <= ~clk;
end
endmodule
